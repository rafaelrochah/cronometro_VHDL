LIBRARY ieee;
USE ieee.std_logic_1164.all;

--LIBRARY work;
--USE work.PORTAS.ALL;

ENTITY MUX_4_1 IS
	PORT
	(
		B1 	:	IN	BIT;
		B2 	:	IN	BIT;
		B3	:	IN	BIT;
		B4	:	IN	BIT;
		C1	: 	IN	BIT;
		C2	:	IN	BIT;
		S : OUT BIT
	);
END MUX_4_1;

ARCHITECTURE ESTRUTURAL OF MUX_4_1 IS

COMPONENT PORTA_AND IS
	PORT
	(
		A	:	IN	BIT;
		B 	: 	IN	BIT;
		C	:	IN	BIT;
		S	:	OUT	BIT
	);
END COMPONENT;

COMPONENT PORTA_OR IS
	PORT
	(
		A	:	IN	BIT;
		B	:	IN	BIT;
		C	:	IN	BIT;
		D	:	IN	BIT;
		S	:	OUT BIT
	);
END COMPONENT;

COMPONENT PORTA_NOT IS
	PORT
	(
		A : IN BIT;
		S : OUT BIT
	);
END COMPONENT;

SIGNAL C1_BARRADO,C2_BARRADO, S1, S2, S3, S4: BIT;

BEGIN
	NOT1 : Porta_NOT PORT MAP (C1,C1_BARRADO);
	NOT2 : Porta_NOT PORT MAP (C2,C2_BARRADO);
	
	AND1	: Porta_AND PORT MAP (B1,C1_BARRADO,C2_BARRADO,S1);
	AND2	: Porta_AND PORT MAP (B2,C1_BARRADO,C2,S2);
	AND3	: Porta_AND PORT MAP (B3,C1,C2_BARRADO,S3);
	AND4	: Porta_AND PORT MAP (B4,C1,C2,S4);
	
	OR1		: Porta_OR PORT MAP (S1,S2,S3,S4,S);
END ESTRUTURAL;