LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY Debouncer IS
	PORT(
		CLK			: in STD_LOGIC;
		CHAVE		: in STD_LOGIC;
		SAIDA		: out STD_LOGIC
		);
END Debouncer;

ARCHITECTURE MISTA OF Debouncer IS

SIGNAL SHIFT_REG : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

	SAIDA <= NOT(SHIFT_REG(0) OR SHIFT_REG(1) OR SHIFT_REG(2) OR SHIFT_REG(3));

	Shift_Register : PROCESS(CLK, CHAVE)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			SHIFT_REG(0) <= CHAVE;
			SHIFT_REG(3 DOWNTO 1) <= SHIFT_REG(2 DOWNTO 0);
		END IF;
	END PROCESS;

END;